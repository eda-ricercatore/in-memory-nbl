*	This is written by Zhiyang
