*	This is written by Zhiyang Ong to model an inverter
*		using 5 um MOSFET devices.
*
*	References:
*		+ \cite[\S8.2, pp. 109; \S8.3.1, pp. 112; \S8.6, pp. 115; \S12.2, pp. 157]{Keiter2019}.
*		+ This specific netlist is from + \cite[\S8.6, pp. 115]{Keiter2019}.


* Subcircuit representation for an inverter,
*	using a 5 um semiconductor manufacturing process technology
.subckt inverter Vin1 Vout Vvdd Vgnd
MN1 VOUT IN 0 0 CD4012_NMOS L=5u W=175u
MP1 VOUT IN VDD VDD CD4012_PMOS L=5u W=270u
.ends


* Schematic of the transistor-level circuit containing an inverter.
VDDdev VDD 0 5V
RIN IN 1 1K
VIN1 1 0 5V PULSE (5V 0V 1.5us 5ns 5ns 1.5us 3us)
R1 VOUT 0 10K
C2 VOUT 0 0.1p
.MODEL cd4012_pmos PMOS
.MODEL cd4012_nmos NMOS
inv in vout Vvdd 0 inverter


* Continuation Options
.options nonlin continuation=mos

* Perform transient analysis circuit simulation step.
.tran 20ns 30us 0 5ns
.print tran v(vout) v(vin1) v(1)
.options timeint reltol=5e-3 abstol=1e-3


.END
